* EESchema Netlist Version 1.1 (Spice format) creation date: Wed 06 Apr 2016 09:00:07 PM CEST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
C4  Net-_C4-Pad1_ Net-_C1-Pad2_ 6.9pF		
L5  Net-_C1-Pad2_ Net-_C5-Pad1_ 18.7nH		
L4  +3V3 Net-_C4-Pad1_ 18.7nH		
L6  +3V3 Net-_C5-Pad1_ 18.7nH		
RDUMMY1  Net-_L2-Pad2_ GND 1G		
C2  GND Net-_C2-Pad2_ 12.7pF		
L1  Net-_C1-Pad1_ Net-_C2-Pad2_ 15.9nH		
L2  Net-_C2-Pad2_ Net-_L2-Pad2_ 15.9nH		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 100pF		
U2  +3V3 GNDD +3V3 ? Net-_C11-Pad1_ MIC5365-2.85YD5-TR		
C3  +3V3 GNDD 1uF		
C11  Net-_C11-Pad1_ GNDD 1uF		
C12  Net-_C11-Pad1_ GNDD 10nF		
C13  Net-_C13-Pad1_ GND 470pF		
C14  Net-_C13-Pad1_ Net-_C14-Pad2_ 6.8nF		
R4  Net-_C14-Pad2_ GND 6.2k		
R5  VTUNE Net-_C13-Pad1_ 13k		
C15  VTUNE GND 220pF		
U3  GNDD GNDD Net-_U1-Pad16_ Net-_C11-Pad1_ XTC7005		
P2  ? ? +3V3 +3V3 GNDD GNDD ? GNDD ? ? ? ? ? ? ? ? ? ? ? ? ? ? PC104		
C5  Net-_C5-Pad1_ GND 6.9pF		
L3  GND GNDD 1mH		

.end
