** ngspice test file for modem filters

.include temp.cir

V1 +3V3 GND 3.3V
I1 NetC4Pad1 GND DC 0 pulse(0mA 11mA      0ns 0.01ns 0.01ns 1.1574ns 2.3148ns)
I2 NetC5Pad1 GND DC 0 pulse(0mA 11mA 1.1574ns 0.01ns 0.01ns 1.1574ns 2.3148ns)
RLOAD NetL2Pad2 temp 50
VLOAD temp GND 0
.tran 0.01ns 2000ns
*the print below shows us 1.29 mW
*print mean( i(vload)^2*50)
.print tran i(vload) v(NetC1Pad1)
.end

